module full_adder (
    input a,
    input b,
    input cin,
    output sum,
    output cout
);
    // Logika Full Adder menggunakan operator bitwise
    assign sum = a ^ b ^ cin;
    assign cout = (a & b) | (b & cin) | (a & cin);

endmodule